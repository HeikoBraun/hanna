LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY design_1 IS
    PORT(
        a: IN    unsigned(3 DOWNTO 0);
        z:   OUT unsigned(3 DOWNTO 0)
    );
END ENTITY design_1;

ARCHITECTURE rtl OF design_1 IS
BEGIN

    z <= a + 2;

END ARCHITECTURE rtl;
