
PACKAGE package_22_pkg IS
    
END PACKAGE package_22_pkg;

