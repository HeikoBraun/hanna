LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ARCHITECTURE rtl OF design_1 IS
BEGIN

    z <= a + 1;
    
END ARCHITECTURE rtl;
