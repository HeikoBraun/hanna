

PACKAGE BODY package_20_pkg IS
    
END PACKAGE BODY package_20_pkg;
