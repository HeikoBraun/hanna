LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ENTITY design_1 IS
    PORT(
        a: IN    std_ulogic;
        z:   OUT std_ulogic
    );
END ENTITY design_1;

