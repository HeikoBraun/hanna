
use work.package_21_pkg.all;
use work.package_22_pkg.all;

PACKAGE package_20_pkg IS
    
END PACKAGE package_20_pkg;
