
PACKAGE package_1_pkg IS
    
END PACKAGE package_1_pkg;
