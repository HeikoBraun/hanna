
CONFIGURATION cfg_design_2 OF design_1 IS
    FOR structure
    END FOR;
END CONFIGURATION cfg_design_2;
