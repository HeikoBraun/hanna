LIBRARY IEEE;
USE ieee.std_logic_1164.all;

LIBRARY lib_2;
USE lib_2.package_20.ALL;
USE lib_2.package_22.ALL;

ARCHITECTURE rtl OF design_1 IS
BEGIN

    z <= a + 1;
    
END ARCHITECTURE rtl;
