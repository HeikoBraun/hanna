module mem_2(a,b,c)
endmodule