
PACKAGE package_21_pkg IS
    
END PACKAGE package_21_pkg;

PACKAGE BODY package_21_pkg IS
    
END PACKAGE BODY package_21_pkg;