
CONFIGURATION cfg_design_1 OF design_1 IS
    FOR rtl
    END FOR;
END CONFIGURATION cfg_design_1;
