module mem_1(a,b,c)
endmodule